library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
use work.timers.all;

entity timer_controller is
    port(inp_switch:in std_logic_vector(2 downto 0);
    reset,clock_50, clock_1:in std_logic;
    out_LED: out std_logic_vector(3 downto 0));
end timer_controller;

architecture behav of timer_controller is

type state is (RST,timer1,timer2,timer3) ;
signal y_present,y_next : state;
signal timer_inp:std_logic_vector(1 downto 0);
component timer_ckt is
    port ( clock_1, clock_50, reset : in std_logic;
    LED : out std_logic_vector(3 downto 0);
    timer_inp : in std_logic_vector(1 downto 0));
end component timer_ckt;

begin
clock_proc:process(clock_50,reset)
begin
    if(clock_50='1' and clock_50' event) then
        if(reset='1') then
            y_present<= RST;
        else
            y_present <= y_next;
        end if;
    end if;
end process ;

state_transition:process(inp_switch,y_present)
begin
    case y_present is
            
            when y_present =>  
            if(inp_switch = 001) then    
                y_next<= timer1;
            elsif(inp_switch= 010) then    
                y_next<= timer2;
            elsif(inp_switch= 100) then    
                y_next<= timer3;
            else 
              y_next <= y_present;
            
            
            end if;
	end case;
end process;
Process(y_present)
begin 
    case y_present is 
        when RST=>
        timer_input := 00;
        when timer1=>
        timer_input := 01;
        when timer2=>
        timer_input := 10;
        when timer3=>
        timer_input := 11;
    end case;
end process;

timer_ckt_1 : timer_ckt port map(clock_1,clock_50,reset,out_LED,timer_input);

end architecture behav;